`include "CPU_wrapper.sv"
`include "AXI/AXI.sv"
`include "SRAM_wrapper.sv"
`include "ROM_wrapper.sv"
`include "DRAM_wrapper.sv"
`include "SC_wrapper.sv"
`include "WDT_wrapper.sv"
//_sdf -version 2.1 -context verilog -load_delay net
module top(
  input clk,
  input clk2,
  input rst,
  input rst2,
  input sensor_ready,
  input [31:0] sensor_out,
  output sensor_en,
  input [31:0] ROM_out,
  input [31:0] DRAM_Q,
  output ROM_read,
  output ROM_enable,
  output [11:0] ROM_address,
  output DRAM_CSn,
  output [3:0] DRAM_WEn,
  output DRAM_RASn,
  output DRAM_CASn,
  output [10:0] DRAM_A,
  output [31:0] DRAM_D,
  input DRAM_valid
);

logic [3:0] AWID_M1;
logic [31:0] AWADDR_M1;
logic [3:0] AWLEN_M1;
logic [2:0] AWSIZE_M1;
logic [1:0] AWBURST_M1;
logic AWVALID_M1;
logic AWREADY_M1;
logic [31:0] WDATA_M1;
logic [3:0] WSTRB_M1;
logic WLAST_M1;
logic WVALID_M1;
logic WREADY_M1;
logic [3:0] BID_M1;
logic [1:0] BRESP_M1;
logic BVALID_M1;
logic BREADY_M1;
////////////////////////////
logic [3:0] ARID_M0,ARID_M1;
logic [31:0] ARADDR_M0,ARADDR_M1;
logic [3:0] ARLEN_M0,ARLEN_M1;
logic [2:0] ARSIZE_M0,ARSIZE_M1;
logic [1:0] ARBURST_M0,ARBURST_M1;
logic ARVALID_M0,ARVALID_M1;
logic ARREADY_M0,ARREADY_M1;
logic [3:0] RID_M0,RID_M1;
logic [31:0] RDATA_M0,RDATA_M1;
logic [1:0] RRESP_M0,RRESP_M1;
logic RLAST_M0,RLAST_M1;
logic RVALID_M0,RVALID_M1;
logic RREADY_M0,RREADY_M1;
///////////////////////////
logic [7:0] AWID_S1,AWID_S2,AWID_S4,AWID_S3,AWID_S5;
logic [31:0] AWADDR_S1,AWADDR_S2,AWADDR_S4,AWADDR_S3,AWADDR_S5;
logic [3:0] AWLEN_S1,AWLEN_S2,AWLEN_S4,AWLEN_S3,AWLEN_S5;
logic [2:0] AWSIZE_S1,AWSIZE_S2,AWSIZE_S4,AWSIZE_S3,AWSIZE_S5;
logic [1:0] AWBURST_S1,AWBURST_S2,AWBURST_S4,AWBURST_S3,AWBURST_S5;
logic AWVALID_S1,AWVALID_S2,AWVALID_S4,AWVALID_S3,AWVALID_S5;
logic AWREADY_S1,AWREADY_S2,AWREADY_S4,AWREADY_S3,AWREADY_S5;
	//WRITE DATA0
logic [31:0] WDATA_S1,WDATA_S2,WDATA_S3,WDATA_S4,WDATA_S5;
logic [3:0] WSTRB_S1,WSTRB_S2,WSTRB_S3,WSTRB_S4,WSTRB_S5;
logic WLAST_S1,WLAST_S2,WLAST_S3,WLAST_S4,WLAST_S5;
logic WVALID_S1,WVALID_S2,WVALID_S3,WVALID_S4,WVALID_S5;
logic WREADY_S1,WREADY_S2,WREADY_S3,WREADY_S4,WREADY_S5;
	//WRITE RESPONSE0
logic [7:0] BID_S1,BID_S2,BID_S3,BID_S4,BID_S5;
logic [1:0] BRESP_S1,BRESP_S2,BRESP_S3,BRESP_S4,BRESP_S5;
logic BVALID_S1,BVALID_S2,BVALID_S3,BVALID_S4,BVALID_S5;
logic BREADY_S1,BREADY_S2,BREADY_S3,BREADY_S4,BREADY_S5;
//READ ADDRESS0
logic [7:0] ARID_S0,ARID_S1,ARID_S2,ARID_S3,ARID_S4,ARID_S5;
logic [31:0] ARADDR_S0,ARADDR_S1,ARADDR_S2,ARADDR_S3,ARADDR_S4,ARADDR_S5;
logic [3:0] ARLEN_S0,ARLEN_S1,ARLEN_S2,ARLEN_S3,ARLEN_S4,ARLEN_S5;
logic [2:0] ARSIZE_S0,ARSIZE_S1,ARSIZE_S2,ARSIZE_S3,ARSIZE_S4,ARSIZE_S5;
logic [1:0] ARBURST_S0,ARBURST_S1,ARBURST_S2,ARBURST_S3,ARBURST_S4,ARBURST_S5;
logic ARVALID_S0,ARVALID_S1,ARVALID_S2,ARVALID_S3,ARVALID_S4,ARVALID_S5;
logic ARREADY_S0,ARREADY_S1,ARREADY_S2,ARREADY_S3,ARREADY_S4,ARREADY_S5;
	//READ DATA0
logic [7:0] RID_S0,RID_S1,RID_S2,RID_S3,RID_S4,RID_S5;
logic [31:0] RDATA_S0,RDATA_S1,RDATA_S2,RDATA_S3,RDATA_S4,RDATA_S5;
logic [1:0] RRESP_S0,RRESP_S1,RRESP_S2,RRESP_S3,RRESP_S4,RRESP_S5;
logic RLAST_S0,RLAST_S1,RLAST_S2,RLAST_S3,RLAST_S4,RLAST_S5;
logic RVALID_S0,RVALID_S1,RVALID_S2,RVALID_S3,RVALID_S4,RVALID_S5;
logic RREADY_S0,RREADY_S1,RREADY_S2,RREADY_S3,RREADY_S4,RREADY_S5;
logic core_interrupt,WDT_interrupt;

CPU_wrapper CP1(
  .clk(clk),.rst(rst),
  //WRITE ADDRESS
	.AWID_M1(AWID_M1),.AWADDR_M1(AWADDR_M1),.AWLEN_M1(AWLEN_M1),.AWSIZE_M1(AWSIZE_M1),
  .AWBURST_M1(AWBURST_M1),.AWVALID_M1(AWVALID_M1),.AWREADY_M1(AWREADY_M1),
	//WRITE DATA
	.WDATA_M1(WDATA_M1),.WSTRB_M1(WSTRB_M1),.WLAST_M1(WLAST_M1),.WVALID_M1(WVALID_M1),.WREADY_M1(WREADY_M1),
	//WRITE RESPONSE
	.BID_M1(BID_M1),.BRESP_M1(BRESP_M1),.BVALID_M1(BVALID_M1),.BREADY_M1(BREADY_M1),

	//READ ADDRESS0 for IM
	.ARID_M0(ARID_M0),.ARADDR_M0(ARADDR_M0),.ARLEN_M0(ARLEN_M0),.ARSIZE_M0(ARSIZE_M0),
  .ARBURST_M0(ARBURST_M0),.ARVALID_M0(ARVALID_M0),.ARREADY_M0(ARREADY_M0),
	//READ DATA0
	.RID_M0(RID_M0),.RDATA_M0(RDATA_M0),.RRESP_M0(RRESP_M0),.RLAST_M0(RLAST_M0),
  .RVALID_M0(RVALID_M0),.RREADY_M0(RREADY_M0),

	//READ ADDRESS1 for DM
	.ARID_M1(ARID_M1),.ARADDR_M1(ARADDR_M1),.ARLEN_M1(ARLEN_M1),.ARSIZE_M1(ARSIZE_M1),
  .ARBURST_M1(ARBURST_M1),.ARVALID_M1(ARVALID_M1),.ARREADY_M1(ARREADY_M1),
	//READ DATA1
	.RID_M1(RID_M1),.RDATA_M1(RDATA_M1),.RRESP_M1(RRESP_M1),.RLAST_M1(RLAST_M1),
  .RVALID_M1(RVALID_M1),.RREADY_M1(RREADY_M1),
  .intr_ex(core_interrupt),
  .intr_tr(WDT_interrupt)
);

AXI AXI1(
  .ACLK(clk),.ARESETn(~rst),
	//SLAVE INTERFACE FOR MASTERS
	//READ ADDRESS0
	.ARID_M0(ARID_M0),.ARADDR_M0(ARADDR_M0),.ARLEN_M0(ARLEN_M0),.ARSIZE_M0(ARSIZE_M0),
  .ARBURST_M0(ARBURST_M0),.ARVALID_M0(ARVALID_M0),.ARREADY_M0(ARREADY_M0),
	//READ DATA0
	.RID_M0(RID_M0),.RDATA_M0(RDATA_M0),.RRESP_M0(RRESP_M0),.RLAST_M0(RLAST_M0),
  .RVALID_M0(RVALID_M0),.RREADY_M0(RREADY_M0),

  .AWID_M1(AWID_M1),.AWADDR_M1(AWADDR_M1),.AWLEN_M1(AWLEN_M1),.AWSIZE_M1(AWSIZE_M1),
  .AWBURST_M1(AWBURST_M1),.AWVALID_M1(AWVALID_M1),.AWREADY_M1(AWREADY_M1),
	//WRITE DATA
	.WDATA_M1(WDATA_M1),.WSTRB_M1(WSTRB_M1),.WLAST_M1(WLAST_M1),.WVALID_M1(WVALID_M1),.WREADY_M1(WREADY_M1),
	//WRITE RESPONSE
	.BID_M1(BID_M1),.BRESP_M1(BRESP_M1),.BVALID_M1(BVALID_M1),.BREADY_M1(BREADY_M1),
	//READ ADDRESS1
	.ARID_M1(ARID_M1),.ARADDR_M1(ARADDR_M1),.ARLEN_M1(ARLEN_M1),.ARSIZE_M1(ARSIZE_M1),
  .ARBURST_M1(ARBURST_M1),.ARVALID_M1(ARVALID_M1),.ARREADY_M1(ARREADY_M1),
	//READ DATA1
	.RID_M1(RID_M1),.RDATA_M1(RDATA_M1),.RRESP_M1(RRESP_M1),.RLAST_M1(RLAST_M1),
  .RVALID_M1(RVALID_M1),.RREADY_M1(RREADY_M1),

	//MASTER INTERFACE FOR SLAVES
	//READ ADDRESS0
	.ARID_S0(ARID_S0),.ARADDR_S0(ARADDR_S0),.ARLEN_S0(ARLEN_S0),.ARSIZE_S0(ARSIZE_S0),
  .ARBURST_S0(ARBURST_S0),.ARVALID_S0(ARVALID_S0),.ARREADY_S0(ARREADY_S0),
	//READ DATA0
  .RID_S0(RID_S0),.RDATA_S0(RDATA_S0),.RRESP_S0(RRESP_S0),.RLAST_S0(RLAST_S0),
  .RVALID_S0(RVALID_S0),.RREADY_S0(RREADY_S0),

	//WRITE ADDRESS1
	.AWID_S1(AWID_S1),.AWADDR_S1(AWADDR_S1),.AWLEN_S1(AWLEN_S1),.AWSIZE_S1(AWSIZE_S1),
  .AWBURST_S1(AWBURST_S1),.AWVALID_S1(AWVALID_S1),.AWREADY_S1(AWREADY_S1),
	//WRITE DATA1
	.WDATA_S1(WDATA_S1),.WSTRB_S1(WSTRB_S1),.WLAST_S1(WLAST_S1),.WVALID_S1(WVALID_S1),.WREADY_S1(WREADY_S1),
	//WRITE RESPONSE1
  .BID_S1(BID_S1),.BRESP_S1(BRESP_S1),.BVALID_S1(BVALID_S1),.BREADY_S1(BREADY_S1),
  //READ ADDRESS1
	.ARID_S1(ARID_S1),.ARADDR_S1(ARADDR_S1),.ARLEN_S1(ARLEN_S1),.ARSIZE_S1(ARSIZE_S1),
  .ARBURST_S1(ARBURST_S1),.ARVALID_S1(ARVALID_S1),.ARREADY_S1(ARREADY_S1),
	//READ DATA1
  .RID_S1(RID_S1),.RDATA_S1(RDATA_S1),.RRESP_S1(RRESP_S1),.RLAST_S1(RLAST_S1),
  .RVALID_S1(RVALID_S1),.RREADY_S1(RREADY_S1),

  //WRITE ADDRESS2
  .AWID_S2(AWID_S2),.AWADDR_S2(AWADDR_S2),.AWLEN_S2(AWLEN_S2),.AWSIZE_S2(AWSIZE_S2),
  .AWBURST_S2(AWBURST_S2),.AWVALID_S2(AWVALID_S2),.AWREADY_S2(AWREADY_S2),
  //WRITE DATA2
  .WDATA_S2(WDATA_S2),.WSTRB_S2(WSTRB_S2),.WLAST_S2(WLAST_S2),.WVALID_S2(WVALID_S2),.WREADY_S2(WREADY_S2),
  //WRITE RESPONSE2
  .BID_S2(BID_S2),.BRESP_S2(BRESP_S2),.BVALID_S2(BVALID_S2),.BREADY_S2(BREADY_S2),
  //READ ADDRESS2
  .ARID_S2(ARID_S2),.ARADDR_S2(ARADDR_S2),.ARLEN_S2(ARLEN_S2),.ARSIZE_S2(ARSIZE_S2),
  .ARBURST_S2(ARBURST_S2),.ARVALID_S2(ARVALID_S2),.ARREADY_S2(ARREADY_S2),
  //READ DATA2
  .RID_S2(RID_S2),.RDATA_S2(RDATA_S2),.RRESP_S2(RRESP_S2),.RLAST_S2(RLAST_S2),
  .RVALID_S2(RVALID_S2),.RREADY_S2(RREADY_S2),

  //WRITE ADDRESS3
  .AWID_S3(AWID_S3),.AWADDR_S3(AWADDR_S3),.AWLEN_S3(AWLEN_S3),.AWSIZE_S3(AWSIZE_S3),
  .AWBURST_S3(AWBURST_S3),.AWVALID_S3(AWVALID_S3),.AWREADY_S3(AWREADY_S3),
  //WRITE DATA3
  .WDATA_S3(WDATA_S3),.WSTRB_S3(WSTRB_S3),.WLAST_S3(WLAST_S3),.WVALID_S3(WVALID_S3),.WREADY_S3(WREADY_S3),
  //WRITE RESPONSE3
  .BID_S3(BID_S3),.BRESP_S3(BRESP_S3),.BVALID_S3(BVALID_S3),.BREADY_S3(BREADY_S3),
  //READ ADDRESS3
  .ARID_S3(ARID_S3),.ARADDR_S3(ARADDR_S3),.ARLEN_S3(ARLEN_S3),.ARSIZE_S3(ARSIZE_S3),
  .ARBURST_S3(ARBURST_S3),.ARVALID_S3(ARVALID_S3),.ARREADY_S3(ARREADY_S3),
  //READ DATA3
  .RID_S3(RID_S3),.RDATA_S3(RDATA_S3),.RRESP_S3(RRESP_S3),.RLAST_S3(RLAST_S3),
  .RVALID_S3(RVALID_S3),.RREADY_S3(RREADY_S3),

  //WRITE ADDRESS4
  .AWID_S4(AWID_S4),.AWADDR_S4(AWADDR_S4),.AWLEN_S4(AWLEN_S4),.AWSIZE_S4(AWSIZE_S4),
  .AWBURST_S4(AWBURST_S4),.AWVALID_S4(AWVALID_S4),.AWREADY_S4(AWREADY_S4),
  //WRITE DATA4
  .WDATA_S4(WDATA_S4),.WSTRB_S4(WSTRB_S4),.WLAST_S4(WLAST_S4),.WVALID_S4(WVALID_S4),.WREADY_S4(WREADY_S4),
  //WRITE RESPONSE4
  .BID_S4(BID_S4),.BRESP_S4(BRESP_S4),.BVALID_S4(BVALID_S4),.BREADY_S4(BREADY_S4),
  //READ ADDRESS4
  .ARID_S4(ARID_S4),.ARADDR_S4(ARADDR_S4),.ARLEN_S4(ARLEN_S4),.ARSIZE_S4(ARSIZE_S4),
  .ARBURST_S4(ARBURST_S4),.ARVALID_S4(ARVALID_S4),.ARREADY_S4(ARREADY_S4),
  //READ DATA4
  .RID_S4(RID_S4),.RDATA_S4(RDATA_S4),.RRESP_S4(RRESP_S4),.RLAST_S4(RLAST_S4),
  .RVALID_S4(RVALID_S4),.RREADY_S4(RREADY_S4),
  
  //WRITE ADDRESS5
  .AWID_S5(AWID_S5),.AWADDR_S5(AWADDR_S5),.AWLEN_S5(AWLEN_S5),.AWSIZE_S5(AWSIZE_S5),
  .AWBURST_S5(AWBURST_S5),.AWVALID_S5(AWVALID_S5),.AWREADY_S5(AWREADY_S5),
  //WRITE DATA5
  .WDATA_S5(WDATA_S5),.WSTRB_S5(WSTRB_S5),.WLAST_S5(WLAST_S5),.WVALID_S5(WVALID_S5),.WREADY_S5(WREADY_S5),
  //WRITE RESPONSE5
  .BID_S5(BID_S5),.BRESP_S5(BRESP_S5),.BVALID_S5(BVALID_S5),.BREADY_S5(BREADY_S5),
  //READ ADDRESS5
  .ARID_S5(ARID_S5),.ARADDR_S5(ARADDR_S5),.ARLEN_S5(ARLEN_S5),.ARSIZE_S5(ARSIZE_S5),
  .ARBURST_S5(ARBURST_S5),.ARVALID_S5(ARVALID_S5),.ARREADY_S5(ARREADY_S5),
  //READ DATA5
  .RID_S5(RID_S5),.RDATA_S5(RDATA_S5),.RRESP_S5(RRESP_S5),.RLAST_S5(RLAST_S5),
  .RVALID_S5(RVALID_S5),.RREADY_S5(RREADY_S5)
);

SRAM_wrapper DM1(
  .CK(clk),.arst(~rst),
  .AWID_S0(AWID_S2),
  .AWADDR_S0(AWADDR_S2),
  .AWLEN_S0(AWLEN_S2),
  .AWSIZE_S0(AWSIZE_S2),
  .AWBURST_S0(AWBURST_S2),
  .AWVALID_S0(AWVALID_S2),
  .AWREADY_S0(AWREADY_S2),
	//WRITE DATA0
  .WDATA_S0(WDATA_S2),
  .WSTRB_S0(WSTRB_S2),
  .WLAST_S0(WLAST_S2),
  .WVALID_S0(WVALID_S2),
  .WREADY_S0(WREADY_S2),
	//WRITE RESPONSE0
  .BID_S0(BID_S2),
  .BRESP_S0(BRESP_S2),
  .BVALID_S0(BVALID_S2),
  .BREADY_S0(BREADY_S2),
  //READ ADDRESS0
  .ARID_S0(ARID_S2),
  .ARADDR_S0(ARADDR_S2),
  .ARLEN_S0(ARLEN_S2),
  .ARSIZE_S0(ARSIZE_S2),
  .ARBURST_S0(ARBURST_S2),
  .ARVALID_S0(ARVALID_S2),
  .ARREADY_S0(ARREADY_S2),
	//READ DATA0
  .RID_S0(RID_S2),
  .RDATA_S0(RDATA_S2),
  .RRESP_S0(RRESP_S2),
  .RLAST_S0(RLAST_S2),
  .RVALID_S0(RVALID_S2),
  .RREADY_S0(RREADY_S2)
);
SRAM_wrapper IM1(
  .CK(clk),.arst(~rst),
  .AWID_S0(AWID_S1),
  .AWADDR_S0(AWADDR_S1),
  .AWLEN_S0(AWLEN_S1),
  .AWSIZE_S0(AWSIZE_S1),
  .AWBURST_S0(AWBURST_S1),
  .AWVALID_S0(AWVALID_S1),
  .AWREADY_S0(AWREADY_S1),
	//WRITE DATA0
  .WDATA_S0(WDATA_S1),
  .WSTRB_S0(WSTRB_S1),
  .WLAST_S0(WLAST_S1),
  .WVALID_S0(WVALID_S1),
  .WREADY_S0(WREADY_S1),
	//WRITE RESPONSE0
  .BID_S0(BID_S1),
  .BRESP_S0(BRESP_S1),
  .BVALID_S0(BVALID_S1),
  .BREADY_S0(BREADY_S1),
  //READ ADDRESS0
  .ARID_S0(ARID_S1),
  .ARADDR_S0(ARADDR_S1),
  .ARLEN_S0(ARLEN_S1),
  .ARSIZE_S0(ARSIZE_S1),
  .ARBURST_S0(ARBURST_S1),
  .ARVALID_S0(ARVALID_S1),
  .ARREADY_S0(ARREADY_S1),
	//READ DATA0
  .RID_S0(RID_S1),
  .RDATA_S0(RDATA_S1),
  .RRESP_S0(RRESP_S1),
  .RLAST_S0(RLAST_S1),
  .RVALID_S0(RVALID_S1),
  .RREADY_S0(RREADY_S1)
);

ROM_wrapper RO1(
  .CK(clk),
  .arst(~rst),
  //READ ADDRESS0
  .ARID_S0(ARID_S0),
  .ARADDR_S0(ARADDR_S0),
  .ARLEN_S0(ARLEN_S0),
  .ARSIZE_S0(ARSIZE_S0),
  .ARBURST_S0(ARBURST_S0),
  .ARVALID_S0(ARVALID_S0),
  .ARREADY_S0(ARREADY_S0),

  .RID_S0(RID_S0),
  .RDATA_S0(RDATA_S0),
  .RRESP_S0(RRESP_S0),
  .RLAST_S0(RLAST_S0),
  .RVALID_S0(RVALID_S0),
  .RREADY_S0(RREADY_S0),
  .ROM_out(ROM_out),
  .ROM_read(ROM_read),
  .ROM_enable(ROM_enable),
  .ROM_address(ROM_address)
);/*
DRAM_wrapper DRA1(
  .CK(clk),
  .arst(~rst),
  //WRITE ADDRESS0
  .AWID_S0(AWID_S4),
  .AWADDR_S0(AWADDR_S4),
  .AWLEN_S0(AWLEN_S4),
  .AWSIZE_S0(AWSIZE_S4),
  .AWBURST_S0(AWBURST_S4),
  .AWVALID_S0(AWVALID_S4),
  .AWREADY_S0(AWREADY_S4),
	//WRITE DATA0
  .WDATA_S0(WDATA_S4),
  .WSTRB_S0(WSTRB_S4),
  .WLAST_S0(WLAST_S4),
  .WVALID_S0(WVALID_S4),
  .WREADY_S0(WREADY_S4),
	//WRITE RESPONSE0
  .BID_S0(BID_S4),
  .BRESP_S0(BRESP_S4),
  .BVALID_S0(BVALID_S4),
  .BREADY_S0(BREADY_S4),
  //READ ADDRESS0
  .ARID_S0(ARID_S4),
  .ARADDR_S0(ARADDR_S4),
  .ARLEN_S0(ARLEN_S4),
  .ARSIZE_S0(ARSIZE_S4),
  .ARBURST_S0(ARBURST_S4),
  .ARVALID_S0(ARVALID_S4),
  .ARREADY_S0(ARREADY_S4),

  .RID_S0(RID_S4),
  .RDATA_S0(RDATA_S4),
  .RRESP_S0(RRESP_S4),
  .RLAST_S0(RLAST_S4),
  .RVALID_S0(RVALID_S4),
  .RREADY_S0(RREADY_S4),
  .DRAM_Q(DRAM_Q),
  .DRAM_CSn(DRAM_CSn),
  .DRAM_WEn(DRAM_WEn),
  .DRAM_RASn(DRAM_RASn),
  .DRAM_CASn(DRAM_CASn),
  .DRAM_A(DRAM_A),
  .DRAM_D(DRAM_D),
	.DRAM_valid(DRAM_valid)
);*/
DRAM_wrapper DRA1(
  .ACLK(clk),
  .ARESETn(~rst),
  //WRITE ADDRESS0
  .AWID(AWID_S5),
  .AWADDR(AWADDR_S5),
  .AWLEN(AWLEN_S5),
  .AWSIZE(AWSIZE_S5),
  .AWBURST(AWBURST_S5),
  .AWVALID(AWVALID_S5),
  .AWREADY(AWREADY_S5),
	//WRITE DATA0
  .WDATA(WDATA_S5),
  .WSTRB(WSTRB_S5),
  .WLAST(WLAST_S5),
  .WVALID(WVALID_S5),
  .WREADY(WREADY_S5),
	//WRITE RESPONSE0
  .BID(BID_S5),
  .BRESP(BRESP_S5),
  .BVALID(BVALID_S5),
  .BREADY(BREADY_S5),
  //READ ADDRESS0
  .ARID(ARID_S5),
  .ARADDR(ARADDR_S5),
  .ARLEN(ARLEN_S5),
  .ARSIZE(ARSIZE_S5),
  .ARBURST(ARBURST_S5),
  .ARVALID(ARVALID_S5),
  .ARREADY(ARREADY_S5),

  .RID(RID_S5),
  .RDATA(RDATA_S5),
  .RRESP(RRESP_S5),
  .RLAST(RLAST_S5),
  .RVALID(RVALID_S5),
  .RREADY(RREADY_S5),
  .DRAM_Q(DRAM_Q),
  .DRAM_CSn(DRAM_CSn),
  .DRAM_WEn(DRAM_WEn),
  .DRAM_RASn(DRAM_RASn),
  .DRAM_CASn(DRAM_CASn),
  .DRAM_A(DRAM_A),
  .DRAM_D(DRAM_D),
  .DRAM_valid(DRAM_valid)
);

SC_wrapper SC0(
  .CK(clk),.arst(~rst),
  .AWID_S0(AWID_S3),
  .AWADDR_S0(AWADDR_S3),
  .AWLEN_S0(AWLEN_S3),
  .AWSIZE_S0(AWSIZE_S3),
  .AWBURST_S0(AWBURST_S3),
  .AWVALID_S0(AWVALID_S3),
  .AWREADY_S0(AWREADY_S3),
	//WRITE DATA0
  .WDATA_S0(WDATA_S3),
  .WSTRB_S0(WSTRB_S3),
  .WLAST_S0(WLAST_S3),
  .WVALID_S0(WVALID_S3),
  .WREADY_S0(WREADY_S3),
	//WRITE RESPONSE0
  .BID_S0(BID_S3),
  .BRESP_S0(BRESP_S3),
  .BVALID_S0(BVALID_S3),
  .BREADY_S0(BREADY_S3),
  //READ ADDRESS0
  .ARID_S0(ARID_S3),
  .ARADDR_S0(ARADDR_S3),
  .ARLEN_S0(ARLEN_S3),
  .ARSIZE_S0(ARSIZE_S3),
  .ARBURST_S0(ARBURST_S3),
  .ARVALID_S0(ARVALID_S3),
  .ARREADY_S0(ARREADY_S3),
	//READ DATA0
  .RID_S0(RID_S3),
  .RDATA_S0(RDATA_S3),
  .RRESP_S0(RRESP_S3),
  .RLAST_S0(RLAST_S3),
  .RVALID_S0(RVALID_S3),
  .RREADY_S0(RREADY_S3),
  .SEN_ready(sensor_ready),
  .SEN_out(sensor_out),
  .SEN_en(sensor_en),
  .SCTRL_irupt(core_interrupt)
);

WDT_wrapper WD0(
  .CK(clk),.arst(~rst),
  .clk2(clk2),.rst2(rst2),
  .AWID_S0(AWID_S4),
  .AWADDR_S0(AWADDR_S4),
  .AWLEN_S0(AWLEN_S4),
  .AWSIZE_S0(AWSIZE_S4),
  .AWBURST_S0(AWBURST_S4),
  .AWVALID_S0(AWVALID_S4),
  .AWREADY_S0(AWREADY_S4),
	//WRITE DATA0
  .WDATA_S0(WDATA_S4),
  .WSTRB_S0(WSTRB_S4),
  .WLAST_S0(WLAST_S4),
  .WVALID_S0(WVALID_S4),
  .WREADY_S0(WREADY_S4),
	//WRITE RESPONSE0
  .BID_S0(BID_S4),
  .BRESP_S0(BRESP_S4),
  .BVALID_S0(BVALID_S4),
  .BREADY_S0(BREADY_S4),
  //READ ADDRESS0
  .ARID_S0(ARID_S4),
  .ARADDR_S0(ARADDR_S4),
  .ARLEN_S0(ARLEN_S4),
  .ARSIZE_S0(ARSIZE_S4),
  .ARBURST_S0(ARBURST_S4),
  .ARVALID_S0(ARVALID_S4),
  .ARREADY_S0(ARREADY_S4),
	//READ DATA0
  .RID_S0(RID_S4),
  .RDATA_S0(RDATA_S4),
  .RRESP_S0(RRESP_S4),
  .RLAST_S0(RLAST_S4),
  .RVALID_S0(RVALID_S4),
  .RREADY_S0(RREADY_S4),
  .WTO(WDT_interrupt)
);

endmodule


